module test_tb();




pll_tb pll_tb0 ();


endmodule